LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity dtrigger is
	port(
	clk,rst,D: in STD_LOGIC;
	Q,not_Q: out STD_LOGIC
	);
	end dtrigger;

architecture bhv of dtrigger is
begin
	process(clk,rst)
	begin
	if clk = '1' and clk'event then
		Q <= D;
		not_Q <= not D;
	end if;
	if rst = '1' then
		Q <= '0';
		not_Q <= '1';
	end if;
	end process;
end bhv;
	